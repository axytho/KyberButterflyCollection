`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/28/2023 08:01:01 PM
// Design Name: 
// Module Name: butterfly_dummy
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module butterfly_dummy(

    );
    
Nguyen_butterfly bf1();
butterfly bf2();
butterfly_xing bf3();
butterfly_Ni bf4();
butterfly_Best bf5();
endmodule
